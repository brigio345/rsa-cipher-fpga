library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package CONSTANTS is
 	
 	constant DATA_WIDTH	 : integer := 16;
	constant ADD_WIDTH	 : integer := 8; 
	
end package CONSTANTS;
